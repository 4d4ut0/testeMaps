** Profile: "SCHEMATIC1-Lab4-1"  [ C:\Users\K4tr1n4\Desktop\aqui\lab4-PSpiceFiles\SCHEMATIC1\Lab4-1.sim ] 

** Creating circuit file "Lab4-1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "Z:/OLB_Pspice/ebipolar.lib" 
* From [PSPICE NETLIST] section of C:\Users\K4tr1n4\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
